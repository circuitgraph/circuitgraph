module s27_unrolled_4 (G1_3, G2_4, DFF_1_Q_reg_Q_0, G1_4, G2_2, G3_1, G1_2, G3_0, G0_4, G0_3, G1_0, G3_3, G1_1, G0_2, DFF_2_Q_reg_Q_0, G0_1, G3_4, G3_2, DFF_0_Q_reg_Q_0, G2_0, G2_1, G2_3, G0_0, G17_3, G17_2, DFF_0_Q_reg_D_4, G17_0, DFF_2_Q_reg_D_4, DFF_1_Q_reg_D_4, G17_1, G17_4);
  input G1_3;
  input G2_4;
  input DFF_1_Q_reg_Q_0;
  input G1_4;
  input G2_2;
  input G3_1;
  input G1_2;
  input G3_0;
  input G0_4;
  input G0_3;
  input G1_0;
  input G3_3;
  input G1_1;
  input G0_2;
  input DFF_2_Q_reg_Q_0;
  input G0_1;
  input G3_4;
  input G3_2;
  input DFF_0_Q_reg_Q_0;
  input G2_0;
  input G2_1;
  input G2_3;
  input G0_0;

  output G17_3;
  output G17_2;
  output DFF_0_Q_reg_D_4;
  output G17_0;
  output DFF_2_Q_reg_D_4;
  output DFF_1_Q_reg_D_4;
  output G17_1;
  output G17_4;

  wire G17_3;
  wire unrolled_4_n_8;
  wire unrolled_4_DFF_2_Q_reg_Q;
  wire unrolled_3_DFF_2_Q_reg_D;
  wire unrolled_0_n_12;
  wire DFF_2_Q_reg_D_2;
  wire DFF_1_Q_reg_Q_2;
  wire unrolled_4_G7;
  wire unrolled_3_G6;
  wire unrolled_0_G1;
  wire unrolled_4_n_4;
  wire DFF_0_Q_reg_D_1;
  wire unrolled_3_n_0;
  wire unrolled_4_n_10;
  wire unrolled_0_n_9;
  wire unrolled_4_n_6;
  wire unrolled_1_n_4;
  wire unrolled_4_DFF_0_Q_reg_Q;
  wire unrolled_1_DFF_2_Q_reg_Q;
  wire unrolled_0_DFF_0_Q_reg_D;
  wire unrolled_1_n_5;
  wire unrolled_1_G7;
  wire unrolled_1_n_10;
  wire unrolled_1_DFF_1_Q_reg_Q;
  wire unrolled_0_n_1;
  wire unrolled_0_n_3;
  wire unrolled_0_n_0;
  wire unrolled_0_n_4;
  wire unrolled_3_G7;
  wire unrolled_3_n_2;
  wire unrolled_0_n_6;
  wire unrolled_3_n_6;
  wire DFF_1_Q_reg_D_1;
  wire unrolled_2_n_21;
  wire DFF_0_Q_reg_Q_3;
  wire unrolled_4_G0;
  wire unrolled_0_DFF_2_Q_reg_D;
  wire unrolled_2_G17_driver;
  wire unrolled_4_n_9;
  wire unrolled_4_n_1;
  wire unrolled_0_n_11;
  wire unrolled_4_n_12;
  wire unrolled_1_G2;
  wire unrolled_2_n_6;
  wire unrolled_2_n_5;
  wire unrolled_3_G17_driver;
  wire unrolled_3_G2;
  wire unrolled_2_n_7;
  wire unrolled_4_G5;
  wire unrolled_4_n_2;
  wire unrolled_1_DFF_0_Q_reg_Q;
  wire unrolled_1_n_8;
  wire DFF_2_Q_reg_Q_4;
  wire G17_4;
  wire unrolled_1_n_2;
  wire unrolled_3_DFF_1_Q_reg_D;
  wire DFF_2_Q_reg_D_1;
  wire unrolled_1_n_3;
  wire unrolled_3_DFF_0_Q_reg_D;
  wire unrolled_1_G17_driver;
  wire unrolled_1_G1;
  wire DFF_2_Q_reg_Q_1;
  wire unrolled_1_G3;
  wire DFF_1_Q_reg_D_2;
  wire unrolled_3_G5;
  wire unrolled_4_G17_driver;
  wire unrolled_2_n_0;
  wire unrolled_2_DFF_2_Q_reg_Q;
  wire unrolled_3_n_5;
  wire unrolled_4_n_5;
  wire unrolled_1_n_0;
  wire unrolled_2_G5;
  wire unrolled_3_n_20;
  wire unrolled_2_DFF_2_Q_reg_D;
  wire DFF_2_Q_reg_D_4;
  wire DFF_0_Q_reg_D_0;
  wire DFF_1_Q_reg_D_0;
  wire unrolled_1_DFF_0_Q_reg_D;
  wire DFF_0_Q_reg_D_3;
  wire unrolled_3_n_4;
  wire DFF_2_Q_reg_Q_2;
  wire DFF_1_Q_reg_Q_1;
  wire unrolled_3_DFF_1_Q_reg_Q;
  wire unrolled_0_n_7;
  wire unrolled_2_n_3;
  wire unrolled_2_n_8;
  wire unrolled_0_G7;
  wire unrolled_4_G3;
  wire unrolled_2_n_1;
  wire unrolled_2_DFF_1_Q_reg_Q;
  wire unrolled_2_G2;
  wire unrolled_1_n_20;
  wire unrolled_1_G0;
  wire unrolled_4_n_0;
  wire unrolled_0_n_5;
  wire unrolled_4_G6;
  wire unrolled_0_n_10;
  wire unrolled_1_n_12;
  wire unrolled_3_n_21;
  wire unrolled_1_n_11;
  wire unrolled_3_n_12;
  wire unrolled_0_G17_driver;
  wire unrolled_2_G0;
  wire unrolled_2_G1;
  wire unrolled_4_G1;
  wire DFF_1_Q_reg_D_4;
  wire G17_1;
  wire DFF_1_Q_reg_Q_4;
  wire unrolled_2_n_2;
  wire unrolled_2_n_12;
  wire unrolled_1_n_7;
  wire DFF_2_Q_reg_D_0;
  wire unrolled_2_G7;
  wire unrolled_2_G3;
  wire unrolled_4_n_7;
  wire unrolled_0_G3;
  wire unrolled_2_n_10;
  wire unrolled_0_DFF_0_Q_reg_Q;
  wire unrolled_1_G6;
  wire unrolled_0_DFF_2_Q_reg_Q;
  wire DFF_0_Q_reg_D_4;
  wire G17_0;
  wire DFF_0_Q_reg_D_2;
  wire unrolled_2_n_9;
  wire unrolled_4_n_3;
  wire unrolled_0_G5;
  wire DFF_0_Q_reg_Q_1;
  wire unrolled_1_n_6;
  wire unrolled_0_DFF_1_Q_reg_D;
  wire unrolled_0_G2;
  wire unrolled_0_DFF_1_Q_reg_Q;
  wire unrolled_2_n_20;
  wire unrolled_3_G0;
  wire unrolled_1_DFF_2_Q_reg_D;
  wire DFF_0_Q_reg_Q_2;
  wire unrolled_1_n_1;
  wire unrolled_4_n_20;
  wire DFF_1_Q_reg_D_3;
  wire unrolled_3_n_7;
  wire unrolled_3_n_3;
  wire unrolled_0_G0;
  wire unrolled_4_n_11;
  wire DFF_2_Q_reg_D_3;
  wire unrolled_3_DFF_0_Q_reg_Q;
  wire unrolled_0_n_21;
  wire unrolled_2_n_11;
  wire unrolled_3_n_1;
  wire unrolled_4_DFF_1_Q_reg_Q;
  wire unrolled_3_n_11;
  wire unrolled_0_n_20;
  wire unrolled_2_DFF_0_Q_reg_D;
  wire DFF_0_Q_reg_Q_4;
  wire DFF_1_Q_reg_Q_3;
  wire unrolled_3_n_9;
  wire unrolled_3_DFF_2_Q_reg_Q;
  wire unrolled_3_n_10;
  wire unrolled_2_DFF_1_Q_reg_D;
  wire unrolled_2_DFF_0_Q_reg_Q;
  wire unrolled_1_DFF_1_Q_reg_D;
  wire unrolled_0_n_2;
  wire DFF_2_Q_reg_Q_3;
  wire unrolled_0_n_8;
  wire unrolled_3_G1;
  wire unrolled_4_G2;
  wire unrolled_2_n_4;
  wire unrolled_3_G3;
  wire G17_2;
  wire unrolled_3_n_8;
  wire unrolled_1_G5;
  wire unrolled_4_n_21;
  wire unrolled_1_n_21;
  wire unrolled_2_G6;
  wire unrolled_0_G6;
  wire unrolled_1_n_9;

  buf g_0 (G17_3, unrolled_3_G17_driver);
  nor g_1 (unrolled_4_n_8, unrolled_4_n_4, unrolled_4_G7);
  buf g_2 (unrolled_4_DFF_2_Q_reg_Q, DFF_2_Q_reg_Q_4);
  buf g_3 (unrolled_3_DFF_2_Q_reg_D, unrolled_3_n_6);
  not g_4 (unrolled_0_n_12, unrolled_0_n_11);
  buf g_5 (DFF_2_Q_reg_D_2, unrolled_2_DFF_2_Q_reg_D);
  buf g_6 (DFF_1_Q_reg_Q_2, DFF_1_Q_reg_D_1);
  buf g_7 (unrolled_4_G7, unrolled_4_DFF_2_Q_reg_Q);
  buf g_8 (unrolled_3_G6, unrolled_3_DFF_1_Q_reg_Q);
  buf g_9 (unrolled_0_G1, G1_0);
  nand g_10 (unrolled_4_n_4, unrolled_4_G3, unrolled_4_n_0);
  buf g_11 (DFF_0_Q_reg_D_1, unrolled_1_DFF_0_Q_reg_D);
  not g_12 (unrolled_3_n_0, unrolled_3_G1);
  nor g_13 (unrolled_4_n_10, unrolled_4_n_7, unrolled_4_n_8);
  nand g_14 (unrolled_0_n_9, unrolled_0_n_1, unrolled_0_n_8);
  nor g_15 (unrolled_4_n_6, unrolled_4_G2, unrolled_4_n_3);
  nand g_16 (unrolled_1_n_4, unrolled_1_n_0, unrolled_1_G3);
  buf g_17 (unrolled_4_DFF_0_Q_reg_Q, DFF_0_Q_reg_Q_4);
  buf g_18 (unrolled_1_DFF_2_Q_reg_Q, DFF_2_Q_reg_Q_1);
  buf g_19 (unrolled_0_DFF_0_Q_reg_D, unrolled_0_n_12);
  nand g_20 (unrolled_1_n_5, unrolled_1_n_2, unrolled_1_G6);
  buf g_21 (unrolled_1_G7, unrolled_1_DFF_2_Q_reg_Q);
  nor g_22 (unrolled_1_n_10, unrolled_1_n_7, unrolled_1_n_8);
  buf g_23 (unrolled_1_DFF_1_Q_reg_Q, DFF_1_Q_reg_Q_1);
  not g_24 (unrolled_0_n_1, unrolled_0_G5);
  nor g_25 (unrolled_0_n_3, unrolled_0_G1, unrolled_0_G7);
  not g_26 (unrolled_0_n_0, unrolled_0_G1);
  nand g_27 (unrolled_0_n_4, unrolled_0_n_0, unrolled_0_G3);
  buf g_28 (unrolled_3_G7, unrolled_3_DFF_2_Q_reg_Q);
  not g_29 (unrolled_3_n_2, unrolled_3_G0);
  nor g_30 (unrolled_0_n_6, unrolled_0_n_3, unrolled_0_G2);
  nor g_31 (unrolled_3_n_6, unrolled_3_G2, unrolled_3_n_3);
  buf g_32 (DFF_1_Q_reg_D_1, unrolled_1_DFF_1_Q_reg_D);
  nor g_33 (unrolled_2_n_21, unrolled_2_G5, unrolled_2_n_10);
  buf g_34 (DFF_0_Q_reg_Q_3, DFF_0_Q_reg_D_2);
  buf g_35 (unrolled_4_G0, G0_4);
  buf g_36 (unrolled_0_DFF_2_Q_reg_D, unrolled_0_n_6);
  not g_37 (unrolled_2_G17_driver, unrolled_2_n_20);
  nand g_38 (unrolled_4_n_9, unrolled_4_n_1, unrolled_4_n_8);
  not g_39 (unrolled_4_n_1, unrolled_4_G5);
  nand g_40 (unrolled_0_n_11, unrolled_0_n_9, unrolled_0_G0);
  not g_41 (unrolled_4_n_12, unrolled_4_n_11);
  buf g_42 (unrolled_1_G2, G2_1);
  nor g_43 (unrolled_2_n_6, unrolled_2_G2, unrolled_2_n_3);
  nand g_44 (unrolled_2_n_5, unrolled_2_G6, unrolled_2_n_2);
  not g_45 (unrolled_3_G17_driver, unrolled_3_n_20);
  buf g_46 (unrolled_3_G2, G2_3);
  not g_47 (unrolled_2_n_7, unrolled_2_n_5);
  buf g_48 (unrolled_4_G5, unrolled_4_DFF_0_Q_reg_Q);
  not g_49 (unrolled_4_n_2, unrolled_4_G0);
  buf g_50 (unrolled_1_DFF_0_Q_reg_Q, DFF_0_Q_reg_Q_1);
  nor g_51 (unrolled_1_n_8, unrolled_1_G7, unrolled_1_n_4);
  buf g_52 (DFF_2_Q_reg_Q_4, DFF_2_Q_reg_D_3);
  buf g_53 (G17_4, unrolled_4_G17_driver);
  not g_54 (unrolled_1_n_2, unrolled_1_G0);
  buf g_55 (unrolled_3_DFF_1_Q_reg_D, unrolled_3_n_21);
  buf g_56 (DFF_2_Q_reg_D_1, unrolled_1_DFF_2_Q_reg_D);
  nor g_57 (unrolled_1_n_3, unrolled_1_G7, unrolled_1_G1);
  buf g_58 (unrolled_3_DFF_0_Q_reg_D, unrolled_3_n_12);
  not g_59 (unrolled_1_G17_driver, unrolled_1_n_20);
  buf g_60 (unrolled_1_G1, G1_1);
  buf g_61 (DFF_2_Q_reg_Q_1, DFF_2_Q_reg_D_0);
  buf g_62 (unrolled_1_G3, G3_1);
  buf g_63 (DFF_1_Q_reg_D_2, unrolled_2_DFF_1_Q_reg_D);
  buf g_64 (unrolled_3_G5, unrolled_3_DFF_0_Q_reg_Q);
  not g_65 (unrolled_4_G17_driver, unrolled_4_n_20);
  not g_66 (unrolled_2_n_0, unrolled_2_G1);
  buf g_67 (unrolled_2_DFF_2_Q_reg_Q, DFF_2_Q_reg_Q_2);
  nand g_68 (unrolled_3_n_5, unrolled_3_G6, unrolled_3_n_2);
  nand g_69 (unrolled_4_n_5, unrolled_4_G6, unrolled_4_n_2);
  not g_70 (unrolled_1_n_0, unrolled_1_G1);
  buf g_71 (unrolled_2_G5, unrolled_2_DFF_0_Q_reg_Q);
  nor g_72 (unrolled_3_n_20, unrolled_3_G5, unrolled_3_n_10);
  buf g_73 (unrolled_2_DFF_2_Q_reg_D, unrolled_2_n_6);
  buf g_74 (DFF_2_Q_reg_D_4, unrolled_4_n_6);
  buf g_75 (DFF_0_Q_reg_D_0, unrolled_0_DFF_0_Q_reg_D);
  buf g_76 (DFF_1_Q_reg_D_0, unrolled_0_DFF_1_Q_reg_D);
  buf g_77 (unrolled_1_DFF_0_Q_reg_D, unrolled_1_n_12);
  buf g_78 (DFF_0_Q_reg_D_3, unrolled_3_DFF_0_Q_reg_D);
  nand g_79 (unrolled_3_n_4, unrolled_3_n_0, unrolled_3_G3);
  buf g_80 (DFF_2_Q_reg_Q_2, DFF_2_Q_reg_D_1);
  buf g_81 (DFF_1_Q_reg_Q_1, DFF_1_Q_reg_D_0);
  buf g_82 (unrolled_3_DFF_1_Q_reg_Q, DFF_1_Q_reg_Q_3);
  not g_83 (unrolled_0_n_7, unrolled_0_n_5);
  nor g_84 (unrolled_2_n_3, unrolled_2_G7, unrolled_2_G1);
  nor g_85 (unrolled_2_n_8, unrolled_2_n_4, unrolled_2_G7);
  buf g_86 (unrolled_0_G7, unrolled_0_DFF_2_Q_reg_Q);
  buf g_87 (unrolled_4_G3, G3_4);
  not g_88 (unrolled_2_n_1, unrolled_2_G5);
  buf g_89 (unrolled_2_DFF_1_Q_reg_Q, DFF_1_Q_reg_Q_2);
  buf g_90 (unrolled_2_G2, G2_2);
  nor g_91 (unrolled_1_n_20, unrolled_1_n_10, unrolled_1_G5);
  buf g_92 (unrolled_1_G0, G0_1);
  not g_93 (unrolled_4_n_0, unrolled_4_G1);
  nand g_94 (unrolled_0_n_5, unrolled_0_n_2, unrolled_0_G6);
  buf g_95 (unrolled_4_G6, unrolled_4_DFF_1_Q_reg_Q);
  nor g_96 (unrolled_0_n_10, unrolled_0_n_7, unrolled_0_n_8);
  not g_97 (unrolled_1_n_12, unrolled_1_n_11);
  nor g_98 (unrolled_3_n_21, unrolled_3_G5, unrolled_3_n_10);
  nand g_99 (unrolled_1_n_11, unrolled_1_G0, unrolled_1_n_9);
  not g_100 (unrolled_3_n_12, unrolled_3_n_11);
  not g_101 (unrolled_0_G17_driver, unrolled_0_n_20);
  buf g_102 (unrolled_2_G0, G0_2);
  buf g_103 (unrolled_2_G1, G1_2);
  buf g_104 (unrolled_4_G1, G1_4);
  buf g_105 (DFF_1_Q_reg_D_4, unrolled_4_n_21);
  buf g_106 (G17_1, unrolled_1_G17_driver);
  buf g_107 (DFF_1_Q_reg_Q_4, DFF_1_Q_reg_D_3);
  not g_108 (unrolled_2_n_2, unrolled_2_G0);
  not g_109 (unrolled_2_n_12, unrolled_2_n_11);
  not g_110 (unrolled_1_n_7, unrolled_1_n_5);
  buf g_111 (DFF_2_Q_reg_D_0, unrolled_0_DFF_2_Q_reg_D);
  buf g_112 (unrolled_2_G7, unrolled_2_DFF_2_Q_reg_Q);
  buf g_113 (unrolled_2_G3, G3_2);
  not g_114 (unrolled_4_n_7, unrolled_4_n_5);
  buf g_115 (unrolled_0_G3, G3_0);
  nor g_116 (unrolled_2_n_10, unrolled_2_n_7, unrolled_2_n_8);
  buf g_117 (unrolled_0_DFF_0_Q_reg_Q, DFF_0_Q_reg_Q_0);
  buf g_118 (unrolled_1_G6, unrolled_1_DFF_1_Q_reg_Q);
  buf g_119 (unrolled_0_DFF_2_Q_reg_Q, DFF_2_Q_reg_Q_0);
  buf g_120 (DFF_0_Q_reg_D_4, unrolled_4_n_12);
  buf g_121 (G17_0, unrolled_0_G17_driver);
  buf g_122 (DFF_0_Q_reg_D_2, unrolled_2_DFF_0_Q_reg_D);
  nand g_123 (unrolled_2_n_9, unrolled_2_n_1, unrolled_2_n_8);
  nor g_124 (unrolled_4_n_3, unrolled_4_G7, unrolled_4_G1);
  buf g_125 (unrolled_0_G5, unrolled_0_DFF_0_Q_reg_Q);
  buf g_126 (DFF_0_Q_reg_Q_1, DFF_0_Q_reg_D_0);
  nor g_127 (unrolled_1_n_6, unrolled_1_n_3, unrolled_1_G2);
  buf g_128 (unrolled_0_DFF_1_Q_reg_D, unrolled_0_n_21);
  buf g_129 (unrolled_0_G2, G2_0);
  buf g_130 (unrolled_0_DFF_1_Q_reg_Q, DFF_1_Q_reg_Q_0);
  nor g_131 (unrolled_2_n_20, unrolled_2_G5, unrolled_2_n_10);
  buf g_132 (unrolled_3_G0, G0_3);
  buf g_133 (unrolled_1_DFF_2_Q_reg_D, unrolled_1_n_6);
  buf g_134 (DFF_0_Q_reg_Q_2, DFF_0_Q_reg_D_1);
  not g_135 (unrolled_1_n_1, unrolled_1_G5);
  nor g_136 (unrolled_4_n_20, unrolled_4_G5, unrolled_4_n_10);
  buf g_137 (DFF_1_Q_reg_D_3, unrolled_3_DFF_1_Q_reg_D);
  not g_138 (unrolled_3_n_7, unrolled_3_n_5);
  nor g_139 (unrolled_3_n_3, unrolled_3_G1, unrolled_3_G7);
  buf g_140 (unrolled_0_G0, G0_0);
  nand g_141 (unrolled_4_n_11, unrolled_4_G0, unrolled_4_n_9);
  buf g_142 (DFF_2_Q_reg_D_3, unrolled_3_DFF_2_Q_reg_D);
  buf g_143 (unrolled_3_DFF_0_Q_reg_Q, DFF_0_Q_reg_Q_3);
  nor g_144 (unrolled_0_n_21, unrolled_0_G5, unrolled_0_n_10);
  nand g_145 (unrolled_2_n_11, unrolled_2_n_9, unrolled_2_G0);
  not g_146 (unrolled_3_n_1, unrolled_3_G5);
  buf g_147 (unrolled_4_DFF_1_Q_reg_Q, DFF_1_Q_reg_Q_4);
  nand g_148 (unrolled_3_n_11, unrolled_3_G0, unrolled_3_n_9);
  nor g_149 (unrolled_0_n_20, unrolled_0_G5, unrolled_0_n_10);
  buf g_150 (unrolled_2_DFF_0_Q_reg_D, unrolled_2_n_12);
  buf g_151 (DFF_0_Q_reg_Q_4, DFF_0_Q_reg_D_3);
  buf g_152 (DFF_1_Q_reg_Q_3, DFF_1_Q_reg_D_2);
  nand g_153 (unrolled_3_n_9, unrolled_3_n_1, unrolled_3_n_8);
  buf g_154 (unrolled_3_DFF_2_Q_reg_Q, DFF_2_Q_reg_Q_3);
  nor g_155 (unrolled_3_n_10, unrolled_3_n_7, unrolled_3_n_8);
  buf g_156 (unrolled_2_DFF_1_Q_reg_D, unrolled_2_n_21);
  buf g_157 (unrolled_2_DFF_0_Q_reg_Q, DFF_0_Q_reg_Q_2);
  buf g_158 (unrolled_1_DFF_1_Q_reg_D, unrolled_1_n_21);
  not g_159 (unrolled_0_n_2, unrolled_0_G0);
  buf g_160 (DFF_2_Q_reg_Q_3, DFF_2_Q_reg_D_2);
  nor g_161 (unrolled_0_n_8, unrolled_0_n_4, unrolled_0_G7);
  buf g_162 (unrolled_3_G1, G1_3);
  buf g_163 (unrolled_4_G2, G2_4);
  nand g_164 (unrolled_2_n_4, unrolled_2_n_0, unrolled_2_G3);
  buf g_165 (unrolled_3_G3, G3_3);
  buf g_166 (G17_2, unrolled_2_G17_driver);
  nor g_167 (unrolled_3_n_8, unrolled_3_G7, unrolled_3_n_4);
  buf g_168 (unrolled_1_G5, unrolled_1_DFF_0_Q_reg_Q);
  nor g_169 (unrolled_4_n_21, unrolled_4_G5, unrolled_4_n_10);
  nor g_170 (unrolled_1_n_21, unrolled_1_n_10, unrolled_1_G5);
  buf g_171 (unrolled_2_G6, unrolled_2_DFF_1_Q_reg_Q);
  buf g_172 (unrolled_0_G6, unrolled_0_DFF_1_Q_reg_Q);
  nand g_173 (unrolled_1_n_9, unrolled_1_n_1, unrolled_1_n_8);
endmodule
